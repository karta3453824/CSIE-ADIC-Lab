//------------------------------------------------------//
//- Advanced Digital IC Design                          //
//-                                                     //
//- Exercise: CONVERTER                                 //
//------------------------------------------------------//

`timescale 1ns/1ps

module CONVERTER(in_8_code, out_129_code);

input [7:0] in_8_code;
output reg [128:0] out_129_code;

always@(*) begin
    case(in_8_code)
        8'd0:   out_129_code = 129'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        8'd1:   out_129_code = 129'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001;
        8'd2:   out_129_code = 129'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011;
        8'd3:   out_129_code = 129'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111;
        8'd4:   out_129_code = 129'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111;
        8'd5:   out_129_code = 129'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111;
        8'd6:   out_129_code = 129'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111;
        8'd7:   out_129_code = 129'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111;
        8'd8:   out_129_code = 129'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111;
        8'd9:   out_129_code = 129'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111;
        8'd10:  out_129_code = 129'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111;
        8'd11:  out_129_code = 129'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111;
        8'd12:  out_129_code = 129'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111;
        8'd13:  out_129_code = 129'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111;
        8'd14:  out_129_code = 129'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111;
        8'd15:  out_129_code = 129'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111;
        8'd16:  out_129_code = 129'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111;
        8'd17:  out_129_code = 129'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111;
        8'd18:  out_129_code = 129'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111;
        8'd19:  out_129_code = 129'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111;
        8'd20:  out_129_code = 129'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111;
        8'd21:  out_129_code = 129'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111;
        8'd22:  out_129_code = 129'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111;
        8'd23:  out_129_code = 129'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111;
        8'd24:  out_129_code = 129'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111;
        8'd25:  out_129_code = 129'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111;
        8'd26:  out_129_code = 129'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111;
        8'd27:  out_129_code = 129'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111;
        8'd28:  out_129_code = 129'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111;
        8'd29:  out_129_code = 129'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111;
        8'd30:  out_129_code = 129'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111;
        8'd31:  out_129_code = 129'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111;
        8'd32:  out_129_code = 129'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111;
        8'd33:  out_129_code = 129'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111;
        8'd34:  out_129_code = 129'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111;
        8'd35:  out_129_code = 129'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111;
        8'd36:  out_129_code = 129'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111;
        8'd37:  out_129_code = 129'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111;
        8'd38:  out_129_code = 129'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111;
        8'd39:  out_129_code = 129'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111;
        8'd40:  out_129_code = 129'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111;
        8'd41:  out_129_code = 129'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111;
        8'd42:  out_129_code = 129'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111;
        8'd43:  out_129_code = 129'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111;
        8'd44:  out_129_code = 129'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111;
        8'd45:  out_129_code = 129'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111;
        8'd46:  out_129_code = 129'b000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111;
        8'd47:  out_129_code = 129'b000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111;
        8'd48:  out_129_code = 129'b000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111;
        8'd49:  out_129_code = 129'b000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111;
        8'd50:  out_129_code = 129'b000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111;
        8'd51:  out_129_code = 129'b000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111;
        8'd52:  out_129_code = 129'b000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111;
        8'd53:  out_129_code = 129'b000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111;
        8'd54:  out_129_code = 129'b000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111;
        8'd55:  out_129_code = 129'b000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111;
        8'd56:  out_129_code = 129'b000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111;
        8'd57:  out_129_code = 129'b000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111;
        8'd58:  out_129_code = 129'b000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111;
        8'd59:  out_129_code = 129'b000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111;
        8'd60:  out_129_code = 129'b000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111;
        8'd61:  out_129_code = 129'b000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111;
        8'd62:  out_129_code = 129'b000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111;
        8'd63:  out_129_code = 129'b000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111;
        8'd64:  out_129_code = 129'b000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111;
        8'd65:  out_129_code = 129'b000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111;
        8'd66:  out_129_code = 129'b000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111;
        8'd67:  out_129_code = 129'b000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111;
        8'd68:  out_129_code = 129'b000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111;
        8'd69:  out_129_code = 129'b000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111;
        8'd70:  out_129_code = 129'b000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111;
        8'd71:  out_129_code = 129'b000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111;
        8'd72:  out_129_code = 129'b000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111;
        8'd73:  out_129_code = 129'b000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111;
        8'd74:  out_129_code = 129'b000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111;
        8'd75:  out_129_code = 129'b000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111;
        8'd76:  out_129_code = 129'b000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111;
        8'd77:  out_129_code = 129'b000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111;
        8'd78:  out_129_code = 129'b000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111;
        8'd79:  out_129_code = 129'b000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111;
        8'd80:  out_129_code = 129'b000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111;
        8'd81:  out_129_code = 129'b000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111;
        8'd82:  out_129_code = 129'b000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111;
        8'd83:  out_129_code = 129'b000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111;
        8'd84:  out_129_code = 129'b000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
        8'd85:  out_129_code = 129'b000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
        8'd86:  out_129_code = 129'b000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
        8'd87:  out_129_code = 129'b000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
        8'd88:  out_129_code = 129'b000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
        8'd89:  out_129_code = 129'b000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
        8'd90:  out_129_code = 129'b000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
        8'd91:  out_129_code = 129'b000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
        8'd92:  out_129_code = 129'b000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
        8'd93:  out_129_code = 129'b000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
        8'd94:  out_129_code = 129'b000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
        8'd95:  out_129_code = 129'b000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
        8'd96:  out_129_code = 129'b000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
        8'd97:  out_129_code = 129'b000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
        8'd98:  out_129_code = 129'b000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
        8'd99:  out_129_code = 129'b000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
        8'd100: out_129_code = 129'b000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
        8'd101: out_129_code = 129'b000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
        8'd102: out_129_code = 129'b000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
        8'd103: out_129_code = 129'b000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
        8'd104: out_129_code = 129'b000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
        8'd105: out_129_code = 129'b000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
        8'd106: out_129_code = 129'b000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
        8'd107: out_129_code = 129'b000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
        8'd108: out_129_code = 129'b000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
        8'd109: out_129_code = 129'b000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
        8'd110: out_129_code = 129'b000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
        8'd111: out_129_code = 129'b000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
        8'd112: out_129_code = 129'b000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
        8'd113: out_129_code = 129'b000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
        8'd114: out_129_code = 129'b000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
        8'd115: out_129_code = 129'b000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
        8'd116: out_129_code = 129'b000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
        8'd117: out_129_code = 129'b000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
        8'd118: out_129_code = 129'b000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
        8'd119: out_129_code = 129'b000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
        8'd120: out_129_code = 129'b000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
        8'd121: out_129_code = 129'b000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
        8'd122: out_129_code = 129'b000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
        8'd123: out_129_code = 129'b000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
        8'd124: out_129_code = 129'b000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
        8'd125: out_129_code = 129'b000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
        8'd126: out_129_code = 129'b000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
        8'd127: out_129_code = 129'b001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
    endcase    
end

endmodule

