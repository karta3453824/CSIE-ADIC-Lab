//------------------------------------------------------//
//- Advanced Digital IC Design                          //
//-                                                     //
//- DCO Modeling                                        //
//------------------------------------------------------//
`timescale 1ns/1ps

module DCO(reset, CODE_0, CODE_1, CODE_2, CODE_3, CODE_4, CODE_5, CODE_6, CODE_7, CODE_8, CODE_9, CODE_10, 
CODE_11, CODE_12, CODE_13, CODE_14, CODE_15, CODE_16, CODE_17, CODE_18, CODE_19, CODE_20, 
CODE_21, CODE_22, CODE_23, CODE_24, CODE_25, CODE_26, CODE_27, CODE_28, CODE_29, CODE_30, 
CODE_31, CODE_32, CODE_33, CODE_34, CODE_35, CODE_36, CODE_37, CODE_38, CODE_39, CODE_40, 
CODE_41, CODE_42, CODE_43, CODE_44, CODE_45, CODE_46, CODE_47, CODE_48, CODE_49, CODE_50, 
CODE_51, CODE_52, CODE_53, CODE_54, CODE_55, CODE_56, CODE_57, CODE_58, CODE_59, CODE_60, 
CODE_61, CODE_62, CODE_63, CODE_64, CODE_65, CODE_66, CODE_67, CODE_68, CODE_69, CODE_70, 
CODE_71, CODE_72, CODE_73, CODE_74, CODE_75, CODE_76, CODE_77, CODE_78, CODE_79, CODE_80, 
CODE_81, CODE_82, CODE_83, CODE_84, CODE_85, CODE_86, CODE_87, CODE_88, CODE_89, CODE_90, 
CODE_91, CODE_92, CODE_93, CODE_94, CODE_95, CODE_96, CODE_97, CODE_98, CODE_99, CODE_100, 
CODE_101, CODE_102, CODE_103, CODE_104, CODE_105, CODE_106, CODE_107, CODE_108, CODE_109, CODE_110, 
CODE_111, CODE_112, CODE_113, CODE_114, CODE_115, CODE_116, CODE_117, CODE_118, CODE_119, CODE_120, 
CODE_121, CODE_122, CODE_123, CODE_124, CODE_125, CODE_126, CODE_127, CODE_128, dco_out);

input reset;
input CODE_0, CODE_1, CODE_2, CODE_3, CODE_4, CODE_5; 
input CODE_6, CODE_7, CODE_8, CODE_9, CODE_10, CODE_11; 
input CODE_12, CODE_13, CODE_14, CODE_15, CODE_16, CODE_17; 
input CODE_18, CODE_19, CODE_20, CODE_21, CODE_22, CODE_23; 
input CODE_24, CODE_25, CODE_26, CODE_27, CODE_28, CODE_29; 
input CODE_30, CODE_31, CODE_32, CODE_33, CODE_34, CODE_35; 
input CODE_36, CODE_37, CODE_38, CODE_39, CODE_40, CODE_41; 
input CODE_42, CODE_43, CODE_44, CODE_45, CODE_46, CODE_47; 
input CODE_48, CODE_49, CODE_50, CODE_51, CODE_52, CODE_53; 
input CODE_54, CODE_55, CODE_56, CODE_57, CODE_58, CODE_59; 
input CODE_60, CODE_61, CODE_62, CODE_63, CODE_64, CODE_65; 
input CODE_66, CODE_67, CODE_68, CODE_69, CODE_70, CODE_71; 
input CODE_72, CODE_73, CODE_74, CODE_75, CODE_76, CODE_77; 
input CODE_78, CODE_79, CODE_80, CODE_81, CODE_82, CODE_83; 
input CODE_84, CODE_85, CODE_86, CODE_87, CODE_88, CODE_89; 
input CODE_90, CODE_91, CODE_92, CODE_93, CODE_94, CODE_95; 
input CODE_96, CODE_97, CODE_98, CODE_99, CODE_100, CODE_101; 
input CODE_102, CODE_103, CODE_104, CODE_105, CODE_106, CODE_107; 
input CODE_108, CODE_109, CODE_110, CODE_111, CODE_112, CODE_113; 
input CODE_114, CODE_115, CODE_116, CODE_117, CODE_118, CODE_119; 
input CODE_120, CODE_121, CODE_122, CODE_123, CODE_124, CODE_125; 
input CODE_126, CODE_127, CODE_128; 

output reg dco_out;

wire [128:0] coarse;

initial dco_out = 1'b0;
real period;

assign coarse = {CODE_128, CODE_127, CODE_126, CODE_125, CODE_124, CODE_123, CODE_122, CODE_121, CODE_120, CODE_119, 
                 CODE_118, CODE_117, CODE_116, CODE_115, CODE_114, CODE_113, CODE_112, CODE_111, CODE_110, CODE_109,
                 CODE_108, CODE_107, CODE_106, CODE_105, CODE_104, CODE_103, CODE_102, CODE_101, CODE_100, CODE_99,
                 CODE_98, CODE_97, CODE_96, CODE_95, CODE_94, CODE_93, CODE_92, CODE_91, CODE_90, CODE_89,
                 CODE_88, CODE_87, CODE_86, CODE_85, CODE_84, CODE_83, CODE_82, CODE_81, CODE_80, CODE_79,
                 CODE_78, CODE_77, CODE_76, CODE_75, CODE_74, CODE_73, CODE_72, CODE_71, CODE_70, CODE_69,
                 CODE_68, CODE_67, CODE_66, CODE_65, CODE_64, CODE_63, CODE_62, CODE_61, CODE_60, CODE_59,
                 CODE_58, CODE_57, CODE_56, CODE_55, CODE_54, CODE_53, CODE_52, CODE_51, CODE_50, CODE_49,
                 CODE_48, CODE_47, CODE_46, CODE_45, CODE_44, CODE_43, CODE_42, CODE_41, CODE_40, CODE_39,
                 CODE_38, CODE_37, CODE_36, CODE_35, CODE_34, CODE_33, CODE_32, CODE_31, CODE_30, CODE_29,
                 CODE_28, CODE_27, CODE_26, CODE_25, CODE_24, CODE_23, CODE_22, CODE_21, CODE_20, CODE_19,
                 CODE_18, CODE_17, CODE_16, CODE_15, CODE_14, CODE_13, CODE_12, CODE_11, CODE_10, CODE_9,
                 CODE_8, CODE_7, CODE_6, CODE_5, CODE_4, CODE_3, CODE_2, CODE_1, CODE_0};

always@(coarse) begin
    case(coarse)
        129'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 : period = 7.5023724;
        129'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001 : period = 5.934624;
        129'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011 : period = 4.6849698;
        129'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111 : period = 4.1400365;
        129'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111 : period = 3.6341645;
        129'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111 : period = 3.1758541;
        129'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111 : period = 2.9209431;
        129'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111 : period = 2.6655217;
        129'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111 : period = 2.4314483;
        129'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111 : period = 2.276363;
        129'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111 : period = 2.1284264;
        129'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111 : period = 1.9755881;
        129'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111 : period = 1.8751793;
        129'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111 : period = 1.7763109;
        129'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111 : period = 1.681098;
        129'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111 : period = 1.6034135;
        129'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111 : period = 1.5301781;
        129'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111 : period = 1.4634987;
        129'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111 : period = 1.4076073;
        129'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111 : period = 1.3531038;
        129'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111 : period = 1.3041881;
        129'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111 : period = 1.2569933;
        129'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111 : period = 1.2201676;
        129'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111 : period = 1.1733667;
        129'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111 : period = 1.1398731;
        129'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111 : period = 1.1117672;
        129'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111 : period = 1.0758777;
        129'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111 : period = 1.0466244;
        129'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111 : period = 1.0184122;
        129'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111 : period = 0.9924748287999999;
        129'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111 : period = 0.9691016929999999;
        129'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111 : period = 0.9434166894;
        129'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111 : period = 0.9252610177;
        129'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111 : period = 0.9027659720000001;
        129'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111 : period = 0.8846073083;
        129'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111 : period = 0.8656019933;
        129'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111 : period = 0.8481712465000001;
        129'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111 : period = 0.8334891814000001;
        129'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111 : period = 0.8160777731;
        129'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111 : period = 0.7992793629;
        129'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111 : period = 0.788168313;
        129'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111 : period = 0.7716582374;
        129'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111 : period = 0.7614365610999999;
        129'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111 : period = 0.7491094527000001;
        129'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111 : period = 0.7354087529;
        129'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111 : period = 0.7244972010999999;
        129'b000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111 : period = 0.7136890154000001;
        129'b000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111 : period = 0.7047754472000001;
        129'b000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111 : period = 0.6933357807;
        129'b000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111 : period = 0.6825503374;
        129'b000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111 : period = 0.674934438;
        129'b000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111 : period = 0.6630453833000001;
        129'b000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111 : period = 0.6549516299;
        129'b000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111 : period = 0.6440269308;
        129'b000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111 : period = 0.6374778869000001;
        129'b000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111 : period = 0.6292303729000001;
        129'b000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111 : period = 0.6212726674000001;
        129'b000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111 : period = 0.6168718304;
        129'b000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111 : period = 0.6060505143;
        129'b000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111 : period = 0.5998871888999999;
        129'b000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111 : period = 0.5931309252;
        129'b000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111 : period = 0.5847079166;
        129'b000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111 : period = 0.5799653029999999;
        129'b000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111 : period = 0.5742429213;
        129'b000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111 : period = 0.5673334411;
        129'b000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111 : period = 0.5607352332000001;
        129'b000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111 : period = 0.5557463281;
        129'b000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111 : period = 0.5493562497000001;
        129'b000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111 : period = 0.5459928628999999;
        129'b000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111 : period = 0.5393183944;
        129'b000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111 : period = 0.5347356581;
        129'b000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111 : period = 0.5306545406000001;
        129'b000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111 : period = 0.5255907847;
        129'b000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111 : period = 0.5214111253;
        129'b000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111 : period = 0.5172697538;
        129'b000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111 : period = 0.5120592901;
        129'b000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111 : period = 0.5070293318;
        129'b000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111 : period = 0.5023642411;
        129'b000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111 : period = 0.5005856347000001;
        129'b000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111 : period = 0.4955531317;
        129'b000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111 : period = 0.49285597400000003;
        129'b000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111 : period = 0.4884368609;
        129'b000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111 : period = 0.4833074273;
        129'b000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111 : period = 0.4805484548;
        129'b000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111 : period = 0.4756737395;
        129'b000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111 : period = 0.4723166435;
        129'b000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111 : period = 0.46846470290000003;
        129'b000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111 : period = 0.4669866874;
        129'b000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111 : period = 0.4633685941;
        129'b000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111 : period = 0.458662889;
        129'b000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111 : period = 0.4568291793;
        129'b000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111 : period = 0.4540882249;
        129'b000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111 : period = 0.451947277;
        129'b000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111 : period = 0.4476108219;
        129'b000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111 : period = 0.4446361868;
        129'b000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111 : period = 0.4416839528;
        129'b000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111 : period = 0.4395310046;
        129'b000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111 : period = 0.43676100209999996;
        129'b000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111 : period = 0.43415481240000003;
        129'b000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111 : period = 0.43004045539999997;
        129'b000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111 : period = 0.4285247854;
        129'b000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111 : period = 0.4264192779;
        129'b000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111 : period = 0.4237921743;
        129'b000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111 : period = 0.4207456088;
        129'b000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111 : period = 0.4189253339;
        129'b000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111 : period = 0.4164332627;
        129'b000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111 : period = 0.41476194829999996;
        129'b000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111 : period = 0.4125132784;
        129'b000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111 : period = 0.410728683;
        129'b000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111 : period = 0.4062462041;
        129'b000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111 : period = 0.4057106994;
        129'b000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111 : period = 0.4035036264;
        129'b000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111 : period = 0.4011036145;
        129'b000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111 : period = 0.3977640245;
        129'b000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111 : period = 0.3961986797;
        129'b000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111 : period = 0.3940700366;
        129'b000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111 : period = 0.3936550585;
        129'b000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111 : period = 0.3911152169;
        129'b000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111 : period = 0.38997974399999996;
        129'b000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111 : period = 0.3867958368;
        129'b000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111 : period = 0.38513099110000004;
        129'b000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111 : period = 0.38300807859999997;
        129'b000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111 : period = 0.38151834380000005;
        129'b000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111 : period = 0.3817320434;
        129'b000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111 : period = 0.3791912298;
        129'b000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111 : period = 0.3776432102;
        129'b000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111 : period = 0.37569316579999995;
        129'b001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111 : period = 0.373296195;
    endcase
end

always@(negedge reset)  //DCO work
begin : dco_run
    forever begin : dco_set
        dco_out = ~dco_out;
        #(period/2.0);             
    end
end

always@(posedge reset) begin  //DCO STOP
    begin
        dco_out = 0;
        disable dco_run;  //turn off DCO when reset = 1;
    end
end

endmodule
