//------------------------------------------------------//
//- Advanced Digital IC Design                          //
//-                                                     //
//- Exercise: Design a FSK Modem                        //
//------------------------------------------------------//
`timescale 1ns/1ps
`include "DCO.v"

module FSK_MODEM(RESET, TX_CLK, TX_DATA, FSK_OUT);

  input  RESET, TX_CLK, TX_DATA;
  output FSK_OUT;

  wire [128:0] FSK_KEY;
  reg  [128:0] FSK_reg;

//DCO
DCO DCO(.reset(RESET), 
.CODE_0(FSK_KEY[0]), .CODE_1(FSK_KEY[1]), .CODE_2(FSK_KEY[2]), .CODE_3(FSK_KEY[3]), .CODE_4(FSK_KEY[4]), .CODE_5(FSK_KEY[5]), 
.CODE_6(FSK_KEY[6]), .CODE_7(FSK_KEY[7]), .CODE_8(FSK_KEY[8]), .CODE_9(FSK_KEY[9]), .CODE_10(FSK_KEY[10]), .CODE_11(FSK_KEY[11]), 
.CODE_12(FSK_KEY[12]), .CODE_13(FSK_KEY[13]), .CODE_14(FSK_KEY[14]), .CODE_15(FSK_KEY[15]), .CODE_16(FSK_KEY[16]), .CODE_17(FSK_KEY[17]), 
.CODE_18(FSK_KEY[18]), .CODE_19(FSK_KEY[19]), .CODE_20(FSK_KEY[20]), .CODE_21(FSK_KEY[21]), .CODE_22(FSK_KEY[22]), .CODE_23(FSK_KEY[23]), 
.CODE_24(FSK_KEY[24]), .CODE_25(FSK_KEY[25]), .CODE_26(FSK_KEY[26]), .CODE_27(FSK_KEY[27]), .CODE_28(FSK_KEY[28]), .CODE_29(FSK_KEY[29]), 
.CODE_30(FSK_KEY[30]), .CODE_31(FSK_KEY[31]), .CODE_32(FSK_KEY[32]), .CODE_33(FSK_KEY[33]), .CODE_34(FSK_KEY[34]), .CODE_35(FSK_KEY[35]), 
.CODE_36(FSK_KEY[36]), .CODE_37(FSK_KEY[37]), .CODE_38(FSK_KEY[38]), .CODE_39(FSK_KEY[39]), .CODE_40(FSK_KEY[40]), .CODE_41(FSK_KEY[41]), 
.CODE_42(FSK_KEY[42]), .CODE_43(FSK_KEY[43]), .CODE_44(FSK_KEY[44]), .CODE_45(FSK_KEY[45]), .CODE_46(FSK_KEY[46]), .CODE_47(FSK_KEY[47]), 
.CODE_48(FSK_KEY[48]), .CODE_49(FSK_KEY[49]), .CODE_50(FSK_KEY[50]), .CODE_51(FSK_KEY[51]), .CODE_52(FSK_KEY[52]), .CODE_53(FSK_KEY[53]), 
.CODE_54(FSK_KEY[54]), .CODE_55(FSK_KEY[55]), .CODE_56(FSK_KEY[56]), .CODE_57(FSK_KEY[57]), .CODE_58(FSK_KEY[58]), .CODE_59(FSK_KEY[59]), 
.CODE_60(FSK_KEY[60]), .CODE_61(FSK_KEY[61]), .CODE_62(FSK_KEY[62]), .CODE_63(FSK_KEY[63]), .CODE_64(FSK_KEY[64]), .CODE_65(FSK_KEY[65]), 
.CODE_66(FSK_KEY[66]), .CODE_67(FSK_KEY[67]), .CODE_68(FSK_KEY[68]), .CODE_69(FSK_KEY[69]), .CODE_70(FSK_KEY[70]), .CODE_71(FSK_KEY[71]), 
.CODE_72(FSK_KEY[72]), .CODE_73(FSK_KEY[73]), .CODE_74(FSK_KEY[74]), .CODE_75(FSK_KEY[75]), .CODE_76(FSK_KEY[76]), .CODE_77(FSK_KEY[77]), 
.CODE_78(FSK_KEY[78]), .CODE_79(FSK_KEY[79]), .CODE_80(FSK_KEY[80]), .CODE_81(FSK_KEY[81]), .CODE_82(FSK_KEY[82]), .CODE_83(FSK_KEY[83]), 
.CODE_84(FSK_KEY[84]), .CODE_85(FSK_KEY[85]), .CODE_86(FSK_KEY[86]), .CODE_87(FSK_KEY[87]), .CODE_88(FSK_KEY[88]), .CODE_89(FSK_KEY[89]), 
.CODE_90(FSK_KEY[90]), .CODE_91(FSK_KEY[91]), .CODE_92(FSK_KEY[92]), .CODE_93(FSK_KEY[93]), .CODE_94(FSK_KEY[94]), .CODE_95(FSK_KEY[95]), 
.CODE_96(FSK_KEY[96]), .CODE_97(FSK_KEY[97]), .CODE_98(FSK_KEY[98]), .CODE_99(FSK_KEY[99]), .CODE_100(FSK_KEY[100]), .CODE_101(FSK_KEY[101]), 
.CODE_102(FSK_KEY[102]), .CODE_103(FSK_KEY[103]), .CODE_104(FSK_KEY[104]), .CODE_105(FSK_KEY[105]), .CODE_106(FSK_KEY[106]), .CODE_107(FSK_KEY[107]), 
.CODE_108(FSK_KEY[108]), .CODE_109(FSK_KEY[109]), .CODE_110(FSK_KEY[110]), .CODE_111(FSK_KEY[111]), .CODE_112(FSK_KEY[112]), .CODE_113(FSK_KEY[113]), 
.CODE_114(FSK_KEY[114]), .CODE_115(FSK_KEY[115]), .CODE_116(FSK_KEY[116]), .CODE_117(FSK_KEY[117]), .CODE_118(FSK_KEY[118]), .CODE_119(FSK_KEY[119]), 
.CODE_120(FSK_KEY[120]), .CODE_121(FSK_KEY[121]), .CODE_122(FSK_KEY[122]), .CODE_123(FSK_KEY[123]), .CODE_124(FSK_KEY[124]), .CODE_125(FSK_KEY[125]), 
.CODE_126(FSK_KEY[126]), .CODE_127(FSK_KEY[127]), .CODE_128(FSK_KEY[128]), .FSK_OUT(FSK_OUT));

//FSK Control
always@(posedge TX_CLK or posedge RESET) begin
    if(RESET)
        FSK_reg <= 129'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    else if(TX_DATA)
        FSK_reg <= 129'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
    else
        FSK_reg <= 129'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
end

assign FSK_KEY = FSK_reg;

endmodule
