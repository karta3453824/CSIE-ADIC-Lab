//------------------------------------------------------//
//- Advanced Digital IC Design                          //
//-                                                     //
//- DCO Modeling                                        //
//------------------------------------------------------//

`timescale 1ns/1ps

module DCO(reset, CODE_0, CODE_1, CODE_2, CODE_3, CODE_4, CODE_5, CODE_6, CODE_7, CODE_8, CODE_9, CODE_10, 
CODE_11, CODE_12, CODE_13, CODE_14, CODE_15, CODE_16, CODE_17, CODE_18, CODE_19, CODE_20, 
CODE_21, CODE_22, CODE_23, CODE_24, CODE_25, CODE_26, CODE_27, CODE_28, CODE_29, CODE_30, 
CODE_31, CODE_32, CODE_33, CODE_34, CODE_35, CODE_36, CODE_37, CODE_38, CODE_39, CODE_40, 
CODE_41, CODE_42, CODE_43, CODE_44, CODE_45, CODE_46, CODE_47, CODE_48, CODE_49, CODE_50, 
CODE_51, CODE_52, CODE_53, CODE_54, CODE_55, CODE_56, CODE_57, CODE_58, CODE_59, CODE_60, 
CODE_61, CODE_62, CODE_63, CODE_64, CODE_65, CODE_66, CODE_67, CODE_68, CODE_69, CODE_70, 
CODE_71, CODE_72, CODE_73, CODE_74, CODE_75, CODE_76, CODE_77, CODE_78, CODE_79, CODE_80, 
CODE_81, CODE_82, CODE_83, CODE_84, CODE_85, CODE_86, CODE_87, CODE_88, CODE_89, CODE_90, 
CODE_91, CODE_92, CODE_93, CODE_94, CODE_95, CODE_96, CODE_97, CODE_98, CODE_99, CODE_100, 
CODE_101, CODE_102, CODE_103, CODE_104, CODE_105, CODE_106, CODE_107, CODE_108, CODE_109, CODE_110, 
CODE_111, CODE_112, CODE_113, CODE_114, CODE_115, CODE_116, CODE_117, CODE_118, CODE_119, CODE_120, 
CODE_121, CODE_122, CODE_123, CODE_124, CODE_125, CODE_126, CODE_127, CODE_128, FSK_OUT);

input reset;
input CODE_0, CODE_1, CODE_2, CODE_3, CODE_4, CODE_5; 
input CODE_6, CODE_7, CODE_8, CODE_9, CODE_10, CODE_11; 
input CODE_12, CODE_13, CODE_14, CODE_15, CODE_16, CODE_17; 
input CODE_18, CODE_19, CODE_20, CODE_21, CODE_22, CODE_23; 
input CODE_24, CODE_25, CODE_26, CODE_27, CODE_28, CODE_29; 
input CODE_30, CODE_31, CODE_32, CODE_33, CODE_34, CODE_35; 
input CODE_36, CODE_37, CODE_38, CODE_39, CODE_40, CODE_41; 
input CODE_42, CODE_43, CODE_44, CODE_45, CODE_46, CODE_47; 
input CODE_48, CODE_49, CODE_50, CODE_51, CODE_52, CODE_53; 
input CODE_54, CODE_55, CODE_56, CODE_57, CODE_58, CODE_59; 
input CODE_60, CODE_61, CODE_62, CODE_63, CODE_64, CODE_65; 
input CODE_66, CODE_67, CODE_68, CODE_69, CODE_70, CODE_71; 
input CODE_72, CODE_73, CODE_74, CODE_75, CODE_76, CODE_77; 
input CODE_78, CODE_79, CODE_80, CODE_81, CODE_82, CODE_83; 
input CODE_84, CODE_85, CODE_86, CODE_87, CODE_88, CODE_89; 
input CODE_90, CODE_91, CODE_92, CODE_93, CODE_94, CODE_95; 
input CODE_96, CODE_97, CODE_98, CODE_99, CODE_100, CODE_101; 
input CODE_102, CODE_103, CODE_104, CODE_105, CODE_106, CODE_107; 
input CODE_108, CODE_109, CODE_110, CODE_111, CODE_112, CODE_113; 
input CODE_114, CODE_115, CODE_116, CODE_117, CODE_118, CODE_119; 
input CODE_120, CODE_121, CODE_122, CODE_123, CODE_124, CODE_125; 
input CODE_126, CODE_127, CODE_128; 
output FSK_OUT;

endmodule
